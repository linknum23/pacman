library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.NUMERIC_STD.all;
use work.pacage.all;

entity font_rom is
  port(
    addr  : in  POINT;
    value : in  integer;
    data  : out std_logic
    );
end font_rom;

architecture Behavioral of font_rom is

  type rom_array is array (integer range <>) of std_logic_vector (0 to 7);
  signal rom : rom_array (0 to 223) := (
    --0
    "00000000",
    "00011100",
    "00100110",
    "01100011",
    "01100011",
    "01100011",
    "00110010",
    "00011100",
    --1
    "00000000",
    "00001100",
    "00011100",
    "00001100",
    "00001100",
    "00001100",
    "00001100",
    "00111111",
    --2
    "00000000",
    "00111110",
    "01100011",
    "00000111",
    "00011110",
    "00111100",
    "01110000",
    "01111111",
    --P (3)
    "00000000",
    "01111110",
    "01100011",
    "01100011",
    "01100011",
    "01111110",
    "01100000",
    "01100000",
    --U (4)
    "00000000",
    "01100011",
    "01100011",
    "01100011",
    "01100011",
    "01100011",
    "01100011",
    "00111110",
    --S (5)
    "00000000",
    "00111100",
    "01100110",
    "01100000",
    "00111110",
    "00000011",
    "01100011",
    "00111110",
    --H (6)
    "00000000",
    "01100011",
    "01100011",
    "01100011",
    "01111111",
    "01100011",
    "01100011",
    "01100011",
    --I (7)
    "00000000",
    "00111111",
    "00001100",
    "00001100",
    "00001100",
    "00001100",
    "00001100",
    "00111111",
    --C (8)
    "00000000",
    "00011110",
    "00110011",
    "01100000",
    "01100000",
    "01100000",
    "00110011",
    "00011110",
    --O (9)
    "00000000",
    "00111110",
    "01100011",
    "01100011",
    "01100011",
    "01100011",
    "01100011",
    "00111110",
    --R (10)
    "00000000",
    "01111110",
    "01100011",
    "01100011",
    "01100111",
    "01111100",
    "01101110",
    "01100111",
    --E (11)
    "00000000",
    "01111111",
    "01100000",
    "01100000",
    "01111110",
    "01100000",
    "01100000",
    "01111111",
    --T (12)
    "00000000",
    "00111111",
    "00001100",
    "00001100",
    "00001100",
    "00001100",
    "00001100",
    "00001100",
    --A (13)
    "00000000",
    "00011100",
    "00110110",
    "01100011",
    "01100011",
    "01111111",
    "01100011",
    "01100011",
    --B (14)
    "00000000",
    "01111110",
    "01100011",
    "01100011",
    "01111110",
    "01100011",
    "01100011",
    "01111110",
    --N (15)
    "00000000",
    "01100011",
    "01110011",
    "01111011",
    "01111111",
    "01101111",
    "01100111",
    "01100011",
    --L (16)
    "00000000",
    "00110000",
    "00110000",
    "00110000",
    "00110000",
    "00110000",
    "00110000",
    "00111111",
    --Y (17)
    "00000000",
    "00110011",
    "00110011",
    "00110011",
    "00011110",
    "00001100",
    "00001100",
    "00001100",
    --copyright (18)
    "00111100",
    "01000010",
    "10011001",
    "10100001",
    "10100001",
    "10011001",
    "01000010",
    "00111100",
    --J (19)
    "00000000",
    "00000011",
    "00000011",
    "00000011",
    "00000011",
    "00000011",
    "01100011",
    "00111110",
    --Z (20)
    "00000000",
    "01111111",
    "00000011",
    "00000110",
    "00011100",
    "00110000",
    "01100000",
    "01111111",
    --D (21)
    "00000000",
    "01111100",
    "01100110",
    "01100011",
    "01100011",
    "01100011",
    "01100110",
    "01111100",
    --expl (22)
    "00000000",
    "00001110",
    "00001110",
    "00011100",
    "00011000",
    "00010000",
    "00000000",
    "00100000",
    --G (23)
    "00000000",
    "00011111",
    "00110000",
    "01100000",
    "01100111",
    "01100011",
    "00110011",
    "00011111",
    --M (24)
    "00000000",
    "01100011",
    "01110111",
    "01111111",
    "01111111",
    "01101011",
    "01100011",
    "01100011",
    --V (25)
    "00000000",
    "01100011",
    "01100011",
    "01100011",
    "01100011",
    "00110110",
    "00011100",
    "00001000",
    --dash (26)
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011100",
    "00000000",
    "00000000",
    "00000000",
    --F (27)
    "00000000",
    "01111111",
    "01100000",
    "01100000",
    "01111110",
    "01100000",
    "01100000",
    "01100000"
    );
  signal why, offset  : unsigned(8 downto 0);
  signal ex           : unsigned(4 downto 0);
  signal newy, newoff : unsigned(why'high downto 0);
  signal newx         : unsigned(ex'high downto 0);
begin
  offset <= to_unsigned(value, 5) & "0000";

  why    <= to_unsigned(addr.Y, why'length);
  ex     <= to_unsigned(addr.X, ex'length);
  newoff <= why + offset;
  newy   <= '0' & newoff(newoff'high downto 1);
  newx   <= '0' & ex(ex'high downto 1);
  process(newx, newy, value)

  begin
    data <= '0';
    if value >= 0 then
      data <= rom(to_integer(newy))(to_integer(newx));
    end if;
  end process;

end Behavioral;
