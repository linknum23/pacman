library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.NUMERIC_STD.all;

entity pacman_rom is
  port(
    addr : in  std_logic_vector(7 downto 0);
    data : out std_logic
    );
end pacman_rom;

architecture Behavioral of pacman_rom is

  type rom_array is array (integer range <>) of std_logic_vector (0 to 31);
  constant rom : rom_array (0 to 63) := (
    --0
    "00000000000000011000000000000000",  --1
    "00000000000000111100000000000000",  --2
    "00000000000001111110000000000000",  --3
    "00000000000011111111000000000000",  --4
    "00000000000111111111100000000000",  --5
    "00000000001111111111110000000000",  --6
    "00000000011111111111111000000000",  --7
    "00000000111111111111111100000000",  --8
    "00000001111111111111111110000000",  --9
    "00000011111111111111111111000000",  --10
    "00000111111111111111111111100000",  --11
    "00001111111111111111111111110000",  --12
    "00011111111111111111111111111000",  --13
    "00111111111111111111111111111100",  --14
    "01111111111111111111111111111110",  --15
    "11111111111111111111111111111111",  --16
    "11111111111111111111111111111111",
    "01111111111111111111111111111110",
    "00111111111111111111111111111100",
    "00011111111111111111111111111000",
    "00001111111111111111111111110000",
    "00000111111111111111111111100000",
    "00000011111111111111111111000000",
    "00000001111111111111111110000000",
    "00000000111111111111111100000000",
    "00000000011111111111111000000000",
    "00000000001111111111110000000000",
    "00000000000111111111100000000000",
    "00000000000011111111000000000000",
    "00000000000001111110000000000000",
    "00000000000000111100000000000000",
    "00000000000000011000000000000000",
--1
    "00000000000000011000000000000000",  --1
    "00000000000000111100000000000000",  --2
    "00000000000001111110000000000000",  --3
    "00000000000011111111000000000000",  --4
    "00000000000111111111100000000000",  --5
    "00000000001111111111110000000000",  --6
    "00000000011111111111111000000000",  --7
    "00000000111111111111111100000000",  --8
    "00000001111111111111111000000000",  --9
    "00000011111111111111110000000000",  --10
    "00000111111111111111100000000000",  --11
    "00001111111111111111000000000000",  --12
    "00011111111111111110000000000000",  --13
    "00111111111111111100000000000000",  --14
    "01111111111111111000000000000000",  --15
    "11111111111111110000000000000000",  --16
    "11111111111111110000000000000000",
    "01111111111111111000000000000000",
    "00111111111111111100000000000000",
    "00011111111111111110000000000000",
    "00001111111111111111000000000000",
    "00000111111111111111100000000000",
    "00000011111111111111110000000000",
    "00000001111111111111111000000000",
    "00000000111111111111111100000000",
    "00000000011111111111111000000000",
    "00000000001111111111110000000000",
    "00000000000111111111100000000000",
    "00000000000011111111000000000000",
    "00000000000001111110000000000000",
    "00000000000000111100000000000000",
    "00000000000000011000000000000000",
    );

  signal offset : std_logic_vector(8 downto 0) := (others => '0');
  signal x, y   : integer                      := 0;
begin

  --mult by 16 by shift 4
  offset <= (data_type & "0000") + addr(7 downto 4);
  y      <= to_integer(unsigned(offset));
  x      <= to_integer(unsigned(addr(3 downto 0)));

  process(y, x)
  begin
    data <= '0';
    if y < 63 and y >= 0 then
      data <= rom(y)(x);
    end if;
  end process;

end Behavioral;
