library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.NUMERIC_STD.all;
use work.pacage.all;

entity ghost_rom is
  port(
    addr   : in  POINT;
    dir : in  DIRECTION;
	 mode : in GHOST_DISP_MODE;
	 squiggle : in std_logic;
    data   : out std_logic_vector(1 downto 0)
    );
end ghost_rom;

architecture Behavioral of ghost_rom is

  type rom_array is array (integer range <>) of std_logic_vector (0 to 31);
  constant rom : rom_array (0 to 159) := (

	--eyes up b1
	"00000000000000000000000000000000",
    "00000000000001010101000000000000",
	"00000000111101010101111100000000",
	"00000010111110010110111110000000",
	"00000110101010010110101010010000",
	"00000110101010010110101010010000",
	"00000101101001010101101001010000",
	"00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010101010101010101010101010100",
	 "00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010101010001010101000101010100",
    "00000101000000010100000001010000",
    "00000000000000000000000000000000",
	                                  
	--eyes up b2                      
	"00000000000000000000000000000000",
    "00000000000001010101000000000000",
	"00000000111101010101111100000000",
	"00000010111110010110111110000000",
	"00000110101010010110101010010000",
	"00000110101010010110101010010000",
	"00000101101001010101101001010000",
	"00010101010101010101010101010100",
    "00010101010101010101010101010100",
	 "00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010100010101000001010100010100",
    "00010000000101000001010000000100",
    "00000000000000000000000000000000",
                                      
	--eyes down b1
    "00000000000000000000000000000000",
    "00000000000001010101000000000000",
    "00000000010101010101010100000000",
    "00000001010101010101010101000000",	
	 "00000101101001010101101001010000",
	 "00010110101010010110101010010100",
	 "00010110101010010110101010010100",
	 "00010110111110010110111110010100",
	 "00010101111101010101111101010100",
    "00010101010101010101010101010100", 
	 "00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010101010001010101000101010100",
    "00000101000000010100000001010000",
    "00000000000000000000000000000000",

	--eyes down b2
    "00000000000000000000000000000000",
    "00000000000001010101000000000000",
    "00000000010101010101010100000000",
    "00000001010101010101010101000000",	
	 "00000101101001010101101001010000",
	 "00010110101010010110101010010100",
	 "00010110101010010110101010010100",
	 "00010110111110010110111110010100",
	 "00010101111101010101111101010100",
    "00010101010101010101010101010100", 
	 "00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010100010101000001010100010100",
    "00010000000101000001010000000100",
    "00000000000000000000000000000000",

	--eyes right b1
	"00000000000000000000000000000000",
    "00000000000001010101000000000000",
    "00000000010101010101010100000000",
    "00000001010101010101010101000000",
    "00000101011010010101011010010000",
    "00000101101010100101101010100000",
    "00000101101011110101101011110000",
	 "00010101101011110101101011110100",
	 "00010101011010010101011010010100",
    "00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010101010001010101000101010100",
    "00000101000000010100000001010000",
    "00000000000000000000000000000000",
	
	--eyes right b2
	 "00000000000000000000000000000000",
    "00000000000001010101000000000000",
    "00000000010101010101010100000000",
    "00000001010101010101010101000000",
    "00000101011010010101011010010000",
    "00000101101010100101101010100000",
    "00000101101011110101101011110000",
	 "00010101101011110101101011110100",
	 "00010101011010010101011010010100",
    "00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010100010101000001010100010100",
    "00010000000101000001010000000100",
    "00000000000000000000000000000000",
	--eyes left b1
    "00000000000000000000000000000000",
    "00000000000001010101000000000000",
    "00000000010101010101010100000000",
    "00000001010101010101010101000000",
	 "00000110100101010110100101010000",--
    "00001010101001011010101001010000",
    "00001111101001011111101001010000",
	 "00011111101001011111101001010100",
	 "00010110100101010110100101010100",--
    "00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010101010001010101000101010100",
    "00000101000000010100000001010000",
    "00000000000000000000000000000000",
	--eyes left b2
    "00000000000000000000000000000000",
    "00000000000001010101000000000000",
    "00000000010101010101010100000000",
    "00000001010101010101010101000000",
	 "00000110100101010110100101010000",--
    "00001010101001011010101001010000",
    "00001111101001011111101001010000",
	 "00011111101001011111101001010100",
	 "00010110100101010110100101010100",--
    "00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010101010101010101010101010100",
    "00010100010101000001010100010100",
    "00010000000101000001010000000100",
    "00000000000000000000000000000000",
	 
	--ghost b1
    "00000000000000000000000000000000",
    "00000000000001010101000000000000",
    "00000000010101010101010100000000",
    "00000001010101010101010101000000",
	 "00000101010101010101010101010000",
    "00000101010101010101010101010000",
    "00000101011010010110100101010000",--eyes
	 "00010101011010010110100101010100",
	 "00010101010101010101010101010100", 
    "00010101010101010101010101010100",
    "00010110100101101001011010010100",--squiggle
    "00011001011010010110100101100100",
    "00010101010101010101010101010100",
    "00010101010001010101000101010100",
    "00000101000000010100000001010000",
    "00000000000000000000000000000000",
	--ghost b2
    "00000000000000000000000000000000",
    "00000000000001010101000000000000",
    "00000000010101010101010100000000",
    "00000001010101010101010101000000",
	 "00000101010101010101010101010000",
    "00000101010101010101010101010000", 
    "00000101011010010110100101010000",--eyes
	 "00010101011010010110100101010100",
	 "00010101010101010101010101010100",	    
    "00010101010101010101010101010100",
	 "00010110100101101001011010010100",--squiggle
    "00011001011010010110100101100100",
    "00010101010101010101010101010100",
    "00010100010101000001010100010100",
    "00010000000101000001010000000100",
    "00000000000000000000000000000000"
    );

  signal why : unsigned(8 downto 0);
  signal ex  : unsigned(4 downto 0);
  signal offset : natural range 0 to 511;

begin

  process(dir,squiggle,mode)
  begin
	 if mode /= FRIGHTENED then
		 case dir is
			when UP =>	
				if squiggle = '1' then 
					offset <= 32;
				else
					offset <= 0;
				end if;
			when DOWN =>
				if squiggle = '1' then 
					offset <= 96;
				else
					offset <= 64;
				end if;
			when R =>
				if squiggle = '1' then 
					offset <= 160;
				else
					offset <= 128;
				end if;
			when L =>
				if squiggle = '1' then 
					offset<= 224;
				else
					offset <= 192;
				end if;
			when others =>
				offset <= 192;
		end case;
	 else
		if squiggle = '1' then 
			offset<= 288;
		else
			offset <= 256;
		end if;
	 end if;
  end process;

  why <= to_unsigned(offset + addr.Y, why'length);
  ex  <= to_unsigned(addr.X, ex'length);

  process(why, ex, offset)
    variable newy : unsigned(why'high downto 0);
    variable newx : unsigned(ex'high downto 0);
  begin
    data <= "00";
    newy := '0' & why(why'high downto 1);
    newx := ex(ex'high downto 1) & '0';
    if newy < 255 and newy >= 0 and newx < 32 and newx >= 0 then
      data <= rom(to_integer(newy))(to_integer(newx))&rom(to_integer(newy))(to_integer(newx)+1);
    end if;
  end process;

end Behavioral;