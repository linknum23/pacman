library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity top_level is
	port (
		mclk : in std_logic
	);
end top_level;

architecture Behavioral of top_level is

begin

end Behavioral;

