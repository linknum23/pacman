library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.pacage.all;


entity pacman_manager is
   port(
      clk : std_logic
      
   );
end pacman_manager;

architecture Behavioral of pacman_manager is

begin


end Behavioral;

